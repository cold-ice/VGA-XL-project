LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY COUNTER IS

GENERIC (MAX				: INTEGER;
			DEBUG 			: INTEGER);
PORT(		STROBE  			: IN  STD_LOGIC;
			EN					: IN STD_LOGIC;
			CL					: IN STD_LOGIC;
			COUNT				: OUT INTEGER RANGE 0 TO MAX
);

END COUNTER;

ARCHITECTURE behavioural OF COUNTER IS

SIGNAL COUNT_BUFFER : INTEGER RANGE 0 TO MAX :=DEBUG;

BEGIN

COUNT <= COUNT_BUFFER;

Counter: PROCESS(STROBE, EN, CL)
BEGIN
	IF(EN='1') THEN
		IF(RISING_EDGE(STROBE)) THEN
			IF(COUNT_BUFFER<MAX) THEN
				COUNT_BUFFER <= COUNT_BUFFER+1;
			ELSE
				COUNT_BUFFER<=0;
			END IF;
		END IF;
	ELSIF(CL='1') THEN
		COUNT_BUFFER <= 0;
	--ELSE
			
	END IF;

END PROCESS;

END behavioural;