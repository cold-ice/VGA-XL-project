LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY REGISTER_32BIT IS

PORT(		STROBE  			: IN  STD_LOGIC;
			EN					: IN STD_LOGIC;
			CL					: IN STD_LOGIC;
			COUNT_X			: OUT INTEGER RANGE 0 TO 797
);

END REGISTER_32BIT;

ARCHITECTURE behavioural OF REGISTER_32BIT IS

SIGNAL COUNT_BUFFER : INTEGER RANGE 0 TO 797 :=0;

BEGIN

COUNT_X <= COUNT_BUFFER;

Counter: PROCESS(STROBE, EN, CL)
BEGIN
	IF(EN='1') THEN
		IF(FALLING_EDGE(STROBE)) THEN
			IF(COUNT_BUFFER<797) THEN
				COUNT_BUFFER <= COUNT_BUFFER+1;
			ELSE
				COUNT_BUFFER<=0;
			END IF;
		END IF;
	ELSIF(CL='1') THEN
		COUNT_BUFFER <= 0;
	--ELSE
			
	END IF;

END PROCESS;

END behavioural;